package mailbox_P;
    import transaction_p::*;
    
    mailbox #(virtual interfaceX) vif_mailbox;
    mailbox #(transaction) tr_mailbox;
    
endpackage